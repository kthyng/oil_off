netcdf ini_fennel {

dimensions:
	xi_rho = 252 ;
	xi_u = 251 ;
	xi_v = 252 ;
	eta_rho = 128 ;
	eta_u = 128 ;
	eta_v = 127 ;
	s_rho = 50 ;
    s_w = 51 ;
	tracer = 15 ;
	ocean_time = 1 ; // (0 currently)

variables:
        int spherical ;
                spherical:long_name = "grid type logical switch" ;
                spherical:flag_values = "0, 1" ;
                spherical:flag_meanings = "Cartesian spherical" ;
        int Vtransform ;
                Vtransform:long_name = "vertical terrain-following transformation equation" ;
        int Vstretching ;
                Vstretching:long_name = "vertical terrain-following stretching function" ;
	double theta_s ;
		theta_s:long_name = "S-coordinate surface control parameter" ;
	double theta_b ;
		theta_b:long_name = "S-coordinate bottom control parameter" ;
	double Tcline ;
		Tcline:long_name = "S-coordinate surface/bottom layer width" ;
		Tcline:units = "meter" ;
	double hc ;
		hc:long_name = "S-coordinate parameter, critical depth" ;
		hc:units = "meter" ;
	double s_rho(s_rho) ;
		s_rho:long_name = "S-coordinate at RHO-points" ;
		s_rho:valid_min = -1. ;
		s_rho:valid_max = 0. ;
                s_rho:positive = "up" ;
                s_rho:standard_name = "ocean_s_coordinate_g1" ;
                s_rho:formula_terms = "s: s_rho C: Cs_r eta: zeta depth: h depth_c: hc" ;
	double s_w(s_w) ;
		s_w:long_name = "S-coordinate at W-points" ;
		s_w:valid_min = -1. ;
		s_w:valid_max = 0. ;
                s_w:positive = "up" ;
                s_w:standard_name = "ocean_s_coordinate_g1" ;
                s_w:formula_terms = "s: s_w C: Cs_w eta: zeta depth: h depth_c: hc" ;
	double Cs_r(s_rho) ;
		Cs_r:long_name = "S-coordinate stretching curves at RHO-points" ;
		Cs_r:valid_min = -1. ;
		Cs_r:valid_max = 0. ;
	double Cs_w(s_w) ;
		Cs_w:long_name = "S-coordinate stretching curves at W-points" ;
		Cs_w:valid_min = -1. ;
		Cs_w:valid_max = 0. ;
        double h(eta_rho, xi_rho) ;
                h:long_name = "bathymetry at RHO-points" ;
                h:units = "meter" ;
                h:coordinates = "lon_rho lat_rho" ;
        double ocean_time(ocean_time) ;
                ocean_time:long_name = "time since initialization" ;
                ocean_time:units = "seconds since 1968-05-23 00:00:00 GMT" ;
	float zeta(ocean_time, eta_rho, xi_rho) ;
		zeta:long_name = "free-surface" ;
		zeta:units = "meter" ;
		zeta:time = "ocean_time" ;
	float ubar(ocean_time, eta_u, xi_u) ;
		ubar:long_name = "vertically integrated u-momentum component" ;
		ubar:units = "meter second-1" ;
		ubar:time = "ocean_time" ;
	float vbar(ocean_time, eta_v, xi_v) ;
		vbar:long_name = "vertically integrated v-momentum component" ;
		vbar:units = "meter second-1" ;
		vbar:time = "ocean_time" ;
	float u(ocean_time, s_rho, eta_u, xi_u) ;
		u:long_name = "u-momentum component" ;
		u:units = "meter second-1" ;
		u:time = "ocean_time" ;
	float v(ocean_time, s_rho, eta_v, xi_v) ;
		v:long_name = "v-momentum component" ;
		v:units = "meter second-1" ;
		v:time = "ocean_time" ;
	float temp(ocean_time, s_rho, eta_rho, xi_rho) ;
		temp:long_name = "potential temperature" ;
		temp:units = "Celsius" ;
		temp:time = "ocean_time" ;
	float salt(ocean_time, s_rho, eta_rho, xi_rho) ;
		salt:long_name = "salinity" ;
		salt:time = "ocean_time" ;
	float NO3(ocean_time, s_rho, eta_rho, xi_rho) ;
		NO3:long_name = "nitrate concentration" ;
		NO3:units = "millimole_N03 meter-3" ;
		NO3:time = "ocean_time" ;
	float NH4(ocean_time, s_rho, eta_rho, xi_rho) ;
		NH4:long_name = "ammonium concentration" ;
		NH4:units = "millimole_NH4 meter-3" ;
		NH4:time = "ocean_time" ;
	float chlorophyll(ocean_time, s_rho, eta_rho, xi_rho) ;
		chlorophyll:long_name = "chlorophyll concentration" ;
		chlorophyll:units = "milligrams_chlorophyll meter-3" ;
		chlorophyll:time = "ocean_time" ;
	float phytoplankton(ocean_time, s_rho, eta_rho, xi_rho) ;
		phytoplankton:long_name = "phytoplankton concentration" ;
		phytoplankton:units = "millimole_nitrogen meter-3" ;
		phytoplankton:time = "ocean_time" ;
	float zooplankton(ocean_time, s_rho, eta_rho, xi_rho) ;
		zooplankton:long_name = "zooplankton concentration" ;
		zooplankton:units = "millimole_nitrogen meter-3" ;
		zooplankton:time = "ocean_time" ;
	float LdetritusN(ocean_time, s_rho, eta_rho, xi_rho) ;
		LdetritusN:long_name = "large fraction nitrogen detritus concentration" ;
		LdetritusN:units = "millimole_nitrogen meter-3" ;
		LdetritusN:time = "ocean_time" ;
	float SdetritusN(ocean_time, s_rho, eta_rho, xi_rho) ;
		SdetritusN:long_name = "small fraction nitrogen detritus concentration" ;
		SdetritusN:units = "millimole_nitrogen meter-3" ;
		SdetritusN:time = "ocean_time" ;
	float LdetritusC(ocean_time, s_rho, eta_rho, xi_rho) ;
		LdetritusC:long_name = "large fraction carbon detritus concentration" ;
		LdetritusC:units = "millimole_carbon meter-3" ;
		LdetritusC:time = "ocean_time" ;
	float SdetritusC(ocean_time, s_rho, eta_rho, xi_rho) ;
		SdetritusC:long_name = "small fraction carbon detritus concentration" ;
		SdetritusC:units = "millimole_carbon meter-3" ;
		SdetritusC:time = "ocean_time" ;
	float TIC(ocean_time, s_rho, eta_rho, xi_rho) ;
		TIC:long_name = "total inorganic carbon" ;
		TIC:units = "millimole_carbon meter-3" ;
		TIC:time = "ocean_time" ;
        float Talk(ocean_time, s_rho, eta_rho, xi_rho) ;
                Talk:long_name = "total alkalinity" ;
                Talk:units = "milliequivalents meter-3" ;
                Talk:time = "ocean_time" ;
    float dye_01(ocean_time, s_rho, eta_rho, xi_rho) ;
		dye_01:long_name = "passive tracer" ;
		dye_01:time = "ocean_time" ;
// global attributes:
		:type = "ROMS INITIAL file" ;
		:title = "ROMS Initial fiels for Hydrodynamics and Biology" ;
		:grd_file = "roms_grd.nc" ;

}
